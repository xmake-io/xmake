module main();
  initial
  begin
    $display("hello world!");
    $finish ;
  end
endmodule
